// Our first program will print the classic "hello world"
// message. Here's the full source code.
module main



fn main() {
	println("hello world")
}
