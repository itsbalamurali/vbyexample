// V's _structs_ are typed collections of fields.
// They're useful for grouping data together to form
// records.

module main



// This `person` struct type has `name` and `age` fields.
type person struct {
	name string
	age  int
}

// NewPerson constructs a new person struct with the given name
fn NewPerson(name string) *person {
	// You can safely return a pointer to local variable
	// as a local variable will survive the scope of the function.
	p := person{name: name}
	p.age = 42
	return &p
}

fn main() {

	// This syntax creates a new struct.
	println(person{"Bob", 20})

	// You can name the fields when initializing a struct.
	println(person{name: "Alice", age: 30})

	// Omitted fields will be zero-valued.
	println(person{name: "Fred"})

	// An `&` prefix yields a pointer to the struct.
	println(&person{name: "Ann", age: 40})

	// It's idiomatic to encapsulate new struct creation in constructor fntions
	println(NewPerson("Jon"))

	// Access struct fields with a dot.
	s := person{name: "Sean", age: 50}
	println(s.name)

	// You can also use dots with struct pointers - the
	// pointers are automatically dereferenced.
	sp := &s
	println(sp.age)

	// Structs are mutable.
	sp.age = 51
	println(sp.age)
}
