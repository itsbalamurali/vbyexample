// Branching with `if` and `else` in V is
// straight-forward.

module main



fn main() {

	// Here's a basic example.
	if 7%2 == 0 {
		println("7 is even")
	} else {
		println("7 is odd")
	}

	// You can have an `if` statement without an else.
	if 8%4 == 0 {
		println("8 is divisible by 4")
	}

	// A statement can precede conditionals; any variables
	// declared in this statement are available in all
	// branches.
	if num := 9; num < 0 {
		println(num, "is negative")
	} else if num < 10 {
		println(num, "has 1 digit")
	} else {
		println(num, "has multiple digits")
	}
}

// Note that you don't need parentheses around conditions
// in V, but that the braces are required.
