// We often need our programs to perform operations on
// collections of data, like selecting all items that
// satisfy a given predicate or mapping all items to a new
// collection with a custom function.

// In some languages it's idiomatic to use [generic](http://en.wikipedia.org/wiki/Generic_programming)
// data structures and algorithms. V does not support
// generics; in V it's common to provide collection
// fntions if and when they are specifically needed for
// your program and data types.

// Here are some example collection fntions for slices
// of `strings`. You can use these examples to build your
// own fntions. Note that in some cases it may be
// clearest to just inline the collection-manipulating
// code directly, instead of creating and calling a
// helper function.

module main

import (
	
	"strings"
)

// Index returns the first index of the target string `t`, or
// -1 if no match is found.
fn Index(vs []string, t string) int {
	for i, v := range vs {
		if v == t {
			return i
		}
	}
	return -1
}

// Include returns `true` if the target string t is in the
// slice.
fn Include(vs []string, t string) bool {
	return Index(vs, t) >= 0
}

// Any returns `true` if one of the strings in the slice
// satisfies the predicate `f`.
fn Any(vs []string, f fn(string) bool) bool {
	for _, v := range vs {
		if f(v) {
			return true
		}
	}
	return false
}

// All returns `true` if all of the strings in the slice
// satisfy the predicate `f`.
fn All(vs []string, f fn(string) bool) bool {
	for _, v := range vs {
		if !f(v) {
			return false
		}
	}
	return true
}

// Filter returns a new slice containing all strings in the
// slice that satisfy the predicate `f`.
fn Filter(vs []string, f fn(string) bool) []string {
	vsf := make([]string, 0)
	for _, v := range vs {
		if f(v) {
			vsf = append(vsf, v)
		}
	}
	return vsf
}

// Map returns a new slice containing the results of applying
// the function `f` to each string in the original slice.
fn Map(vs []string, f fn(string) string) []string {
	vsm := make([]string, len(vs))
	for i, v := range vs {
		vsm[i] = f(v)
	}
	return vsm
}

fn main() {

	// Here we try out our various collection fntions.
	var strs = []string{"peach", "apple", "pear", "plum"}

	println(Index(strs, "pear"))

	println(Include(strs, "grape"))

	println(Any(strs, fn(v string) bool {
		return strings.HasPrefix(v, "p")
	}))

	println(All(strs, fn(v string) bool {
		return strings.HasPrefix(v, "p")
	}))

	println(Filter(strs, fn(v string) bool {
		return strings.Contains(v, "e")
	}))

	// The above examples all used anonymous fntions,
	// but you can also use named fntions of the correct
	// type.
	println(Map(strs, strings.ToUpper))

}
